`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:45:23 12/13/2024
// Design Name:   F_Permutation_Dilithium
// Module Name:   C:/Users/fossu/Desktop/SHA3_imp/F_Permutation_Dilithium/F_Permutation_Dilithium_tb.v
// Project Name:  F_Permutation_Dilithium
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: F_Permutation_Dilithium
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module F_Permutation_Dilithium_tb;

	// Inputs
	reg clk;
	reg reset;
	reg [1343:0] in;
	reg in_ready;
	reg squeeze;
	reg [1:0] mode;
	reg sha_hold;

	// Outputs
	wire ack;
	wire [1599:0] out;
	wire out_ready;

	// Instantiate the Unit Under Test (UUT)
	F_Permutation_Dilithium uut (
		.clk(clk), 
		.reset(reset), 
		.in(in), 
		.in_ready(in_ready), 
		.squeeze(squeeze), 
		.mode(mode), 
		.sha_hold(sha_hold), 
		.ack(ack), 
		.out(out), 
		.out_ready(out_ready)
	);

	always begin
		clk = ~clk;
		#5;
	end
	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		in = 0;
		in_ready = 0;
		squeeze = 0;
		mode = 0;
		sha_hold = 0;

		// Wait 100 ns for global reset to finish
		#100;
		reset = 0;
		in = 1600'b1010010111101100101111000110010100110010101000101111010011010111011000000100101011000001100000010110110101101010110111000011010011111101010111101010100111110110101101010101000000011101011010000111000110000101100011101000010000001011101011000000001011010011001000000010000011111000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        mode = 2'b10;
		#10;
		in_ready = 1;
		squeeze = 0;
		// Add stimulus here

	end
      
endmodule

