`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   22:45:23 12/13/2024
// Design Name:   F_Permutation_Dilithium
// Module Name:   C:/Users/fossu/Desktop/SHA3_imp/F_Permutation_Dilithium/F_Permutation_Dilithium_tb.v
// Project Name:  F_Permutation_Dilithium
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: F_Permutation_Dilithium
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module F_Permutation_Dilithium_tb;

	// Inputs
	reg clk;
	reg reset;
	reg [1343:0] in;
	reg in_ready;
	reg squeeze;
	reg [1:0] mode;
	reg sha_hold;

	// Outputs
	wire ack;
	wire [1599:0] out;
	wire out_ready;

	// Instantiate the Unit Under Test (UUT)
	F_Permutation_Dilithium uut (
		.clk(clk), 
		.reset(reset), 
		.in(in), 
		.in_ready(in_ready), 
		.squeeze(squeeze), 
		.mode(mode), 
		.sha_hold(sha_hold), 
		.ack(ack), 
		.out(out), 
		.out_ready(out_ready)
	);

	always begin
		clk = ~clk;
		#5;
	end
	initial begin
		// Initialize Inputs
		clk = 0;
		reset = 1;
		in = 0;
		in_ready = 0;
		squeeze = 0;
		mode = 0;
		sha_hold = 0;

		// Wait 100 ns for global reset to finish
		#100;
		reset = 0;
		// in = 1344'b100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000100000001001100101101000000001101011101000000100001011100011010000110001110000101101011100000001010101011010110111110010101011110101011111100101100001110110101011010110110100000011000001101010010000001101110101100101111010001010100110010100110001111010011011110100101;
		// in = 1344'b101001011110110010111100011001010011001010100010111101001101011101100000010010101100000110000001011011010110101011011100001101001111110101011110101010011111011010110101010100000001110101101000011100011000010110001110100001000000101110101100000000101101001100100000001000001111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001;
		// in = 1344'b110101111111010010100010001100100110010110111100111011001010010100110100110111000110101001101101100000011100000101001010011000000110100000011101010100001011010111110110101010010101111011111101110100110000001010101100000010111000010010001110100001010111000100000000000000000000000000000000000000001111100000100000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000;
		// in = 1344'd0;

		in = 1344'b000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111100000100000001000001101001100000010101011000000101110000100100011101000010101110001011010000001110101010000101101011111011010101001010111101111110100110100110111000110101001101101100000011100000101001010011000001101011111110100101000100011001001100101101111001110110010100101;
        mode = 2'b00;
		#10;
		in_ready = 1;
		squeeze = 0;
		// Add stimulus here

	end

	always @(posedge clk)begin
		if(out_ready)$display("out: %h.", out);
	end
      
endmodule

